CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 3 120 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
3 4 0.500000 0.500000
344 176 457 273
76546066 0
0
6 Title:
5 Name:
0
0
0
11
7 Ground~
168 898 133 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7159 0 0
2
43530.4 0
0
2 +V
167 190 268 0 1 3
0 16
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5812 0 0
2
43530.4 1
0
6 74112~
219 648 352 0 7 32
0 16 15 17 15 16 18 3
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U4B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 4 0
1 U
331 0 0
2
5.89884e-315 0
0
6 74112~
219 495 351 0 7 32
0 16 7 17 7 16 19 6
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U4A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 4 0
1 U
9604 0 0
2
5.89884e-315 5.26354e-315
0
6 74112~
219 333 351 0 7 32
0 16 4 17 4 16 20 5
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 3 0
1 U
7518 0 0
2
5.89884e-315 5.30499e-315
0
6 74112~
219 190 351 0 7 32
0 16 16 17 16 16 21 4
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 3 0
1 U
4832 0 0
2
5.89884e-315 5.32571e-315
0
9 CC 7-Seg~
183 802 152 0 17 19
10 8 9 10 11 12 13 14 22 2
1 1 1 0 0 1 1 2
0
0 0 21104 0
7 AMBERCC
9 -41 58 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
6798 0 0
2
5.89884e-315 5.34643e-315
0
6 74LS48
188 801 323 0 14 29
0 3 6 5 4 23 24 14 13 12
11 10 9 8 25
0
0 0 4848 0
7 74LS248
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3336 0 0
2
5.89884e-315 5.3568e-315
0
9 2-In AND~
219 584 206 0 3 22
0 7 6 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
8370 0 0
2
5.89884e-315 5.36716e-315
0
9 2-In AND~
219 420 204 0 3 22
0 4 5 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3910 0 0
2
5.89884e-315 5.37752e-315
0
7 Pulser~
4 66 317 0 10 12
0 26 27 28 17 0 0 5 5 5
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
316 0 0
2
5.89884e-315 5.38788e-315
0
37
1 0 3 0 0 8336 0 8 0 0 29 5
769 287
738 287
738 411
683 411
683 316
4 0 4 0 0 12416 0 8 0 0 30 5
769 314
755 314
755 428
228 428
228 315
0 3 5 0 0 8320 0 0 8 24 0 5
372 315
372 423
750 423
750 305
769 305
2 0 6 0 0 12416 0 8 0 0 23 5
769 296
744 296
744 417
529 417
529 315
9 1 2 0 0 8320 0 7 1 0 0 4
802 110
802 100
898 100
898 127
0 0 7 0 0 4224 0 0 0 7 19 2
462 204
462 315
3 1 7 0 0 0 0 10 9 0 0 4
441 204
552 204
552 197
560 197
0 1 4 0 0 0 0 0 10 9 0 4
268 316
268 205
396 205
396 195
4 0 4 0 0 0 0 5 0 0 30 3
309 333
268 333
268 315
13 1 8 0 0 8320 0 8 7 0 0 5
833 341
876 341
876 228
781 228
781 188
12 2 9 0 0 8320 0 8 7 0 0 5
833 332
870 332
870 232
787 232
787 188
11 3 10 0 0 8320 0 8 7 0 0 5
833 323
865 323
865 236
793 236
793 188
10 4 11 0 0 8320 0 8 7 0 0 5
833 314
861 314
861 240
799 240
799 188
9 5 12 0 0 8320 0 8 7 0 0 5
833 305
857 305
857 244
805 244
805 188
8 6 13 0 0 16512 0 8 7 0 0 5
833 296
852 296
852 248
811 248
811 188
7 7 14 0 0 16512 0 8 7 0 0 5
833 287
847 287
847 252
817 252
817 188
2 0 15 0 0 4096 0 3 0 0 18 2
624 316
608 316
4 3 15 0 0 8320 0 3 9 0 0 4
624 334
608 334
608 206
605 206
2 4 7 0 0 0 0 4 4 0 0 4
471 315
459 315
459 333
471 333
2 0 16 0 0 4096 0 6 0 0 21 2
166 315
153 315
4 1 16 0 0 8192 0 6 2 0 0 5
166 333
153 333
153 281
190 281
190 277
0 0 16 0 0 4096 0 0 0 27 37 2
244 281
244 372
2 7 6 0 0 0 0 9 4 0 0 4
560 215
540 215
540 315
519 315
2 7 5 0 0 0 0 10 5 0 0 4
396 213
378 213
378 315
357 315
1 0 16 0 0 0 0 5 0 0 27 2
333 288
333 281
1 0 16 0 0 0 0 4 0 0 27 2
495 288
495 281
1 1 16 0 0 8320 0 2 3 0 0 4
190 277
190 281
648 281
648 289
1 1 16 0 0 0 0 2 6 0 0 2
190 277
190 288
7 0 3 0 0 0 0 3 0 0 0 2
672 316
711 316
7 2 4 0 0 0 0 6 5 0 0 2
214 315
309 315
3 0 17 0 0 8192 0 4 0 0 34 3
465 324
451 324
451 396
3 0 17 0 0 0 0 5 0 0 34 3
303 324
288 324
288 396
3 0 17 0 0 0 0 6 0 0 34 3
160 324
145 324
145 396
4 3 17 0 0 12416 0 11 3 0 0 6
96 317
117 317
117 396
603 396
603 325
618 325
5 0 16 0 0 0 0 4 0 0 37 2
495 363
495 372
5 0 16 0 0 0 0 5 0 0 37 2
333 363
333 372
5 5 16 0 0 0 0 6 3 0 0 4
190 363
190 372
648 372
648 364
3
-16 0 0 0 700 255 0 0 0 3 2 1 66
12 Segoe Script
0 0 0 9
9 37 121 79
19 45 110 71
9 BSCPE 1-B
-19 0 0 0 700 255 0 0 0 1 2 1 34
11 Small Fonts
0 0 0 35
214 86 676 116
224 94 665 116
35 BINARY 4-BIT SYNCHRONOUS UP COUNTER
-16 0 0 0 700 255 0 0 0 3 2 1 66
12 Segoe Script
0 0 0 24
9 11 264 53
18 18 254 44
24 TUBAC, CRISTINE DOLOR A.
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
